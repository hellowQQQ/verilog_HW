module top(
		input 		 clk,
		input 		 rstn,
		output [7:0] ledo
		);

	

endmodule